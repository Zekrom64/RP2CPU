module Cpu65EL02DataSeq();

endmodule
